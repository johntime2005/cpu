`timescale 1ns / 1ps

// 此文件内容已被清空，先前的测试平台不再需要。
// 请根据新的测试需求创建或修改测试平台。

module tb_deprecated;
    // 模块内容已移除
endmodule